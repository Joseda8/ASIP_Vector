module vector_reg_bank();




endmodule
